-- MotorPasso_tb.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity MotorPasso_tb is
end entity MotorPasso_tb;

architecture rtl of MotorPasso_tb is
	component MotorPasso is
		port (
			chaves_export : in  std_logic_vector(3 downto 0) := (others => 'X'); -- export
			clk_clk       : in  std_logic                    := 'X';             -- clk
			leds_name     : out std_logic_vector(3 downto 0);                    -- name
			reset_reset_n : in  std_logic                    := 'X'              -- reset_n
		);
	end component MotorPasso;

	component altera_conduit_bfm is
		port (
			sig_export : out std_logic_vector(3 downto 0)   -- export
		);
	end component altera_conduit_bfm;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_conduit_bfm_0002 is
		port (
			clk      : in std_logic                    := 'X';             -- clk
			sig_name : in std_logic_vector(3 downto 0) := (others => 'X'); -- name
			reset    : in std_logic                    := 'X'              -- reset
		);
	end component altera_conduit_bfm_0002;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal motorpasso_inst_clk_bfm_clk_clk           : std_logic;                    -- MotorPasso_inst_clk_bfm:clk -> [MotorPasso_inst:clk_clk, MotorPasso_inst_leds_bfm:clk, MotorPasso_inst_reset_bfm:clk]
	signal motorpasso_inst_chaves_bfm_conduit_export : std_logic_vector(3 downto 0); -- MotorPasso_inst_chaves_bfm:sig_export -> MotorPasso_inst:chaves_export
	signal motorpasso_inst_leds_name                 : std_logic_vector(3 downto 0); -- MotorPasso_inst:leds_name -> MotorPasso_inst_leds_bfm:sig_name
	signal motorpasso_inst_reset_bfm_reset_reset     : std_logic;                    -- MotorPasso_inst_reset_bfm:reset -> MotorPasso_inst:reset_reset_n

begin

	motorpasso_inst : component MotorPasso
		port map (
			chaves_export => motorpasso_inst_chaves_bfm_conduit_export, -- chaves.export
			clk_clk       => motorpasso_inst_clk_bfm_clk_clk,           --    clk.clk
			leds_name     => motorpasso_inst_leds_name,                 --   leds.name
			reset_reset_n => motorpasso_inst_reset_bfm_reset_reset      --  reset.reset_n
		);

	motorpasso_inst_chaves_bfm : component altera_conduit_bfm
		port map (
			sig_export => motorpasso_inst_chaves_bfm_conduit_export  -- conduit.export
		);

	motorpasso_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => motorpasso_inst_clk_bfm_clk_clk  -- clk.clk
		);

	motorpasso_inst_leds_bfm : component altera_conduit_bfm_0002
		port map (
			clk      => motorpasso_inst_clk_bfm_clk_clk, --     clk.clk
			sig_name => motorpasso_inst_leds_name,       -- conduit.name
			reset    => '0'                              -- (terminated)
		);

	motorpasso_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => motorpasso_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => motorpasso_inst_clk_bfm_clk_clk        --   clk.clk
		);

end architecture rtl; -- of MotorPasso_tb
