
module MotorPasso (
	chaves_export,
	clk_clk,
	reset_reset_n,
	phases_phases);	

	input	[3:0]	chaves_export;
	input		clk_clk;
	input		reset_reset_n;
	output	[3:0]	phases_phases;
endmodule
